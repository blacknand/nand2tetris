module not(in, out);
    input in;
    output out;
endmodule